module FFT (clk, rst, s1, l1);
    input clk, rst, data_in;
    output l1;
endmodule