module FFT-H_top (clk, rst, data_in, data_out);
    input clk, rst, data_in;
    output data_out;
endmodule